module divider();

	parameter data_width = 64;


	
endmodule